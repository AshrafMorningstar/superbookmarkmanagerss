-- Created by: Ashraf Morningstar
-- GitHub: https://github.com/AshrafMorningstar

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Hello World does not directly apply, this is a placeholder.
entity hello_world is
end hello_world;

architecture behavioral of hello_world is
begin
end behavioral;