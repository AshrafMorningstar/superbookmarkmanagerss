/*
 Copyright (c) 2026 Ashraf Morningstar
 These are personal recreations of existing projects, developed by Ashraf Morningstar
 for learning and skill development.
 Original project concepts remain the intellectual property of their respective creators.
 Repository: https://github.com/AshrafMorningstar
*/

// Created by: Ashraf Morningstar
// GitHub: https://github.com/AshrafMorningstar

module hello_world;
  initial begin
    $display("Hello, World!");
    $finish;
  end
endmodule