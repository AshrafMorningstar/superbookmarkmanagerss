// Bluespec Test File
// Auto-generated by Ashraf Morningstar
// GitHub: https://github.com/AshrafMorningstar
// Created: 2025-11-13 23:36:45

// This is a test file for Bluespec
// File extension: .bsv
// Auto-generated by Ashraf Morningstar

main_function() {
    print("Hello from Bluespec!");
    return "Hello, World!";
}

// Execute
main_function();