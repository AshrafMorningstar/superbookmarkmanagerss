// Created by: Ashraf Morningstar
// GitHub: https://github.com/AshrafMorningstar

module hello_world;
  initial begin
    $display("Hello, World!");
    $finish;
  end
endmodule